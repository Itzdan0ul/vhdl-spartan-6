----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:26:04 01/06/2023 
-- Design Name: 
-- Module Name:    main_constraints - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity main_constraints is
    Port ( S0 : in  STD_LOGIC;
           S1 : in  STD_LOGIC;
           S2 : in  STD_LOGIC;
           N0 : in  STD_LOGIC;
           N1 : in  STD_LOGIC;
           N2 : in  STD_LOGIC;
           MY : out  STD_LOGIC;
           ME : out  STD_LOGIC;
           EQ : out  STD_LOGIC);
end main_constraints;

architecture Behavioral of main_constraints is

begin


end Behavioral;

